`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.05.2019 13:06:03
// Design Name: 
// Module Name: wcdma_ovsf_generator
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module wcdma_ovsf_generator(
    input aclk,
    input arst,
    input [31:0] axis,
    output [31:0] aixm
    );
endmodule
